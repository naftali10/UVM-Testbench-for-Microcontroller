`include "defines.sv"

package tb_pkg;

  import uvm_pkg::*;
  import definitions::*;

  `include "transaction_class.svh"
  `include "sequence_class.svh"
  `include "sequencer_class.svh"
  `include "driver_class.svh"
  `include "monitor_class.svh"
  `include "agent_class.svh"
  `include "reference_model_class.svh"
  `include "coverage_transaction.sv"
  `include "covergroup_container.sv"
  `include "coverage_analyzer.sv"
  `include "subscriber_class.svh"
  `include "comparator_class.svh"
  `include "scoreboard_class.svh"
  `include "env_class.svh"
  `include "test_class.svh"

endpackage: tb_pkg
