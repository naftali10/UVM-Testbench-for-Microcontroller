`include "defines.sv"		// has to be first
`include "multiplexer.sv"
`include "SHFL.sv"
`include "ALU.sv"
`include "RF.sv"
`include "controller.sv"
`include "reg_out.sv"
`include "reg_EXtoWB.sv"
`include "reg_IDtoEX.sv"
`include "ifc_WB.sv"
`include "ifc_inputs.sv"
`include "Decode.sv"
`include "Execute.sv"
`include "WriteBack.sv"
`include "Top.sv"
`include "ifc_outputs.sv"
`include "Output.sv"
