`include "includes.sv"
